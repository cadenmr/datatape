// Ethernet Data Parser

module ethernet_parse(

	input wire [0:0]	rst,
	input wire [0:0]	clk	// Same as Ethernet clock (125 MHz)

);



endmodule