// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UJamD96X78BrWx8u92nIROC8MCuC3jQq4pMJuvSuWsyzYZ0tvy2ARv0idYXVVuw6FG67NFSj/lEO
go+Bs0AXnzSSTAZIIezTuFyTKWf3fHiwmENnDn7WXScqsBqfJOXbcBd2ZAO/FjYsrWHezoCtBB52
b0D09XkvvRGe+LDO0xq5dfpbkyHqCM2vjGgMWeS9tg0v/PCDRvAQHDVW6RWdGUShl4REOSIOQGCp
laPsQBA85qsBGjZSB2wri0spihFgzdTNY9YGxRm0h2Uh/funvD5WhtdE4XnW+XHhoiFzgJBAUjjQ
GIqk1+EHlPTWn1426Rk4lGPaR09A69B5mP8fDQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5760)
AwMc7XWmCDMNAqsdI9EgSW6ZXPSUDJcMBToce10XoPZAGmRtcdIL7pMBgyxRXNAIwRsXDmKbFeO8
PVf5g43y8WVXvfFGn1yvRbbvUxor/N/mHJ3+Y9zfKJERZ+CZCLtFIejrFEnCfFXh8UiVA8bg7Q+k
FAixHDg43lpbwrXlH565btwU4EVU9JBxoLZ2gwHowsNjEqtdo3MvmvctT06SDp5pQZ86D3C/wP+Q
1wm81mgz7fs8roP32DipY/buXq5ik3L6ItGkXIIBCZOn7CUgvsAepgauI9bCkbGGfXpAyGmXeH79
Zmghjs56Nb0sngWh/rBS/Ew/P5/0YJS1feQN1b9U/vnZSyHhYZT/l1JjSeYm6YpqjMr0YFkGlty3
Fl1MfioyNV7tqZH4UyiHDGQM5hoKrO94tQGjuTLpLB67MnSXmHEqKB6D6vuY8SRg8HwphncUWCVL
SVsW14PydhAEqDCdYxXR3DG6xiFuso4NzEQhw6VvJz//mCrFYUhf+VlUVCI5TsSQ7VkTbJ6eKJew
S73tcx0F/KAOiLFsPLjCHxCvXN7HgLepJpHpY5QvMSp/WbLPIcTIBf6vkBFE5CG/BudTNVheqEPY
KdaW+mYzeOfSKg6NSaVg47xD5v4FNnQNUUgyC9yKYg6j2O1zVurc53w+Dohox+tnaMkMKAv6EYXb
79lsPs7jvJeE7aMlWYgrUPvWYdjZYFQXeJD2AkK+QkKqmFVzUihkeIPZ82zpvHEpSyPB4zUI1O6R
/CAoYDsx+UUTkkWukKL/6UnbeaDKY8/HHjN/3U7Cm3C0gTAZL5uY3Fz2XWVjgKQ0YO/sfT8lGCcX
jGa5t3kt1/2A45zDdnxdxNRTpfD+Cj+08RrQssSsB2Wcxg7M93DAuv8wrprOwYGDhvGibYwW+RcU
WikDh+yHqQCFq5c63xDlIxRbeCU+x86nDPx2ltPjr2logrGcfoN0Qs15N8m9bFKS2uFhMyd3Hu4e
xw+DAXkDAqH5ILjTRKCV30mMLAtj+RibkiYh+kf2vKNj4OrCaZP/Uj24zLcPZZJwzMBxk04FZ16p
KXcRNJCqyA9Mgn3yTMdkfQ7MkZ/0cUhvZ7AH29gjrjOiEJ4BDzwATDZsx7Ui/djjInCqh7vAIidv
sjfqSs4paIMMzcQNsPr+LVa5pHFpgFBRsStL9uNhNqwmQwKNe5UIvjG4KRklzTowYfCRHnMBnytN
QEj2Qmr9M677eLrxbKEUaRrsaXOs849K0RDRLUqV+iucKDjxCQ89j8E5ZOMal0QO7ko4h0oEeozN
1i0DIijoIG5XiMQXg0jW79Z9ImNFWBz7SMAKBS6oXIpRO1bbr3jfZ12NptVKTIPeOM3IM1SIzMEG
khoAXbSZX9a+0fG7mSxUbxTNQ51kJ5a8u7RXVi0yYxy6yjjmoDhAn7dz9kLz3TVOFqTf131WxQwl
V+H/dfIMeEm7DLuXmrMxYCaonCy5PozRnZcrVSl5gWqZxxuVE8UDyYDR4EkVwZUzuCuul8mCU/id
COzKWEbKxQC6bRL90T7Mef/1+hj/5t4cEFC62lWtZ92bMMWMvc1nRAcCsTNCy1rIYamU3vNcL11D
aVlkQbOa0d7BXaRPrPpQ5PIbIpNcX6XhlgIB2gnGTxoGoWP3x1LvnD8B3TvqUGKf2b7Llb1Nxzma
WpcqRb7E2T4W9Uq4XkSyG7I9uobtyoN8e3tPqp+HA7pLEAEXzWUYYdXrvLh7XdBpazsYipGJNteb
twD/Ziub5Deunf5yTibGfLAZmC2p0D+Iblk2fgbCyYAi2OF3YKtXVLJPAbwlRi4vx+bgMrP3px14
x5Qn24c3KCcbVOuqvpSLUf4U5JesaekM3Mmw4GRdOsY+iz5SUfpNWq9yr51Nrjv5hDp4Ll2jDgPs
YLHrLMu1GtUZ3QjJ0OLlpLNv1Wsb8a6z5e+pXFipkmp3PNjHWPPLU3hE1KqJfyTmQ3b2fm0HXBRp
n9LMBzRtyFoFcU1BORiCbh6+/kJ5I5zd9btnnBRVkue01G/X4yjOBUrIiBQBZUCv6qvAHugwuCoF
I7i+j2/P+j37KdVa9Q3xSA4xzt6jJjjlAa3veQw3IUUkZKVg03RJbRARSpv/lLQXpbH7o5deiQlE
V/rO+iPD0FVp86oCRdCToHPLLDDk9Om4DoBNZsyB1EYhdKSlVt2mbotYKEG//7D0QoCSC5CkfTOi
wnTF/0f97nH102IphronGS9JqfCpTlGE2yL6nGO9cMIOzl6SBSfCGXDGN4/D43gh7SEqnbTx/jBt
2F94vMKlaN5c1vBTblcKNoQ2yMOEICtShOAZR8RrwmsJqcbm1VsmKor9RZ1gHlxDSDVAkcxRuV9k
H/krbuyk8QvRWccfuM58DuQVUVPctB/r44toDcbBQahukuMJxIgjD/15pe08p0HuLc2vO3zJaBhY
ZnTlqDf7j0It7m1uqnOvS/1gzJQ7c3So5XpkEZBRxfEOl8IQFZnUk6+JypzxVqgKzI1f+giNP3PX
kCQMD9dQ1khLPN9dLg2rgTnSnjGtAullPg7RIaKN8A3+6UTcYHf3ZQh7qr5n3g3xi3sWXJal0Qdn
HaZHj40KjLR2PlT/taTQ+73YH0dbxeBhf2h8dT40sDfCFkuCM3UrnVPO5yJjfTeIUr/7XDW17r2W
S36HDw5Bra+dFFEGbP5idDFqgE+bNf+KM3mDpTNXt13hxIutchnAJOFu3Lgenv7xwAoHY04Dbz2m
0nUzR4aX0z6WHFAAeyWSb7eMuXgR7h3VTfHxNbDGhnNTyuWXTWmV6I9eFCD4JOYFT0+/hkQiRPmi
rLPHg20cQOFnhlsDWPlyjcPFsyUxWqNnViSOZOO5mW3k+BlkXgEb8wLRRlZXcFtWVVv8xjlKRpAB
qXrkhCeRLW6lI3cVLcmrq7eQh6f2uN5ETydHK9VQL1avpcJPkNrPE+xCVDCTqDWADRrfCz/b/dsE
u24zUFNKGLgLSuvEFBL0KjfSRsk1Z0jg0s4XUaydbjmutOjKTQLSegjDdTtSKikU5clwCK7PEINt
Mm7IeGBOOvQCk/vNaKfgiLfUKKCrCb8M5mNWKbtdUOzhM5z2IvXRJrJPwiai/363zEGA4lUBU4t0
1M6YALzxnNXDE6sIxttl9JDl9d9164x/RLNZ830eEbwUFx3TAWe1aFHMmh9kxZj+v8v/QHeVxa11
VukLyhwx9/h87nUrma+WkzTdCyN5jDdDNk0DLmuyPu+0xEynMBYY5s4sCYnJuJ5WJ0XLtdWSOFXO
Wifu7pt/cHe+S3KUVvkZP5zVAt/SIag6RgxUMMu3osbnmzFJ32GEXQP6QLxYcwcePpy9EkWP8Icv
Zq7ngwywN+9bibGlgqJjZNyNrYLYE5X5KhspM4WsOEGohEQOtgIHW0XjoDKHxtKffnsO/aCnP+z2
5ebCKAh3xll4hJZE0TJbRfz+cg5syimd6l4A2mk3fpSF7Fim78G5LdNmTk0qdWte4eV9rweNyMlj
a/RWgRQu/uLTq5YNhBR387yjJ2aEXT9q9PBkE+KsOLhMvs+TEWTnwkEQJW4a3rg7c+wOI+jbReNX
T0XsSaF0qny+IExG5XJpmkz8BN6VkH/lxruuGt6o0jetvCdhKFyvKf43lj9tQpbnU8vDL9M52rFp
GfD7tuHrx401DYyaADVXVmHfmq/SsnFE0v7L2AZUZYJ/e/RoCgy0DlajmVj8ZhjdJahs6Jx67IzE
yrlIxeLsI5FxITSKRFKL+kIHeQvL+wco3zjLspEfUeSNMsOyRa85yjrVXpA0bKpDcgl4V36xm3gg
9kXM9c1vEBmF4Sb5VhTvPCdoGMWZhyfldJ2pOI54SUdnLoq3G3ItEKexHKDmgFB6JFqovuy3AshH
XkI8whmxFpx9NOE2iaiX7lpR5/hTD4RIEbuPVZYOG9GFyAWr+3o1mrdsDjkDkIXVRsqnBub/ANUS
MyqUntp+xwaGqSiV8hL7AuzFMrAKAFkLJhcLFU+sIIgGZsgJO9YBsw6GguiNP2uv0kImiQ2pbGbt
J7qxrD5dbtAQ2HolirOpkH6hxuPNy7h4s5bwDyPqmPVpEXvkBAmKwtVOBh7qstQ3d53HEB96Laz0
kkHFMjBInyBvNtJXZhs0mRSoo3+rGkzMShtCPGat/fn/ub66jqNLZeBchF7ixINaKm15dqS7l9FB
U9G3iaI7AH+D7FOtt+LcUOTbJLIJ26rCG9zucd0XouABbAl3BDJq9/6tHelw0BW7XfRWdI66ykRR
cgeUfQnDG5W3ABXjBIaPJkhNFcf45o+cxNPi+ElJltS760U2kWiEit87p2ohuRW2Z86Burke4jWg
bJcBV9AKJhJHtayFzzr2sr94pVeD0aAQj/kgNbnqOf1EK4tQSSSGtjHJoFtJ0b9aTGcJtntrMM1g
TK8K9ULdBGLjhTloOG41kvbf/r7jIL0suTJNYApHg+steYfXjcCH+4ZiHyIQIKtSZ1qZcD5mQvdM
sYKODDY5EnDDAfEdO8C59AT2FY2yGK7HsbOmfG418IgVDnuB0SBvMcODTE9wUpUG2gu/jiZtfEM9
rblHuAsBO6rMqPVftnLvXvHyMbj0AHmbO5GqP11wHN2zvoa0qWyd+V2B7UgEf0aQWLp8RzBYABj+
m1YxWScsQiQL/sdc3bmBauINhQ0BUaDPokMTiasGScDzKlZn0PWDUQ9427E0sioG0o8dLGmP5i1m
fMDxllMdZN2jgA4P8U22cBhRCiXe2H5rCpSSOABDwaqRQLkYpW12HJkfKJHIda1r4huxn5vWA/iS
HElz/0hdLO1ZHYxCM9HZv759PnFWzictse+pJ+2juSuU3U57xNZ6OWWXejpsDgyf7ljqA9ohioko
DDdCNRJlVsE1mKtoi1h0U0MIRwq+uKHJe5CbrZ3NhJbsa1bkbmpa6wsx1KrvXPsJnbsocDxh8gqB
sQbTLSRMfJ7PtTn+yaLyNCCtm/TW22Mzyy2S7pyUnF7edHT1TcRAGysyifniLXykCNQdb52tFSk1
8+OlZ7vHrbAKilv8bE4x8hstIF8U9M25k/4ST+yagdfwRW3rWVNXtqf7ue9rxmu1VuDxAOmw6MFR
Lzk7yvyaSgZXXoO0Igiqs9rRFqzSk2LzPm+f7v5Vv95CPExQx2ml8sROJIFFmfHwhSQugtg1KMqn
DyJgKt5UQxKALNwOZqm8EmcFuT8t8zR9Iz6u85uu2ieohLIb+FIqzineRMVQRQF1aoS9ErjBPyU6
w7Y8yqx359Cy1gB5GwOFQwOQQIdOiOKORw4d6b9QvtP5jG7mZOGmqa+BpoLDu2Rh1RrACu/bLR93
bV54mIndt1lTBpo2eTcBG/YfOrRJbkit/aMZQU3rH4AOtEfaniwknXToIDh0ulAA/bN6KrEWIFQ8
Dzbhj4w8Q5JBneCHo8aTcEjCV77lo44pcr6QUnRQtXexCJflhShjOhPT+wS5/rLclo0ELlBfz62J
ofMqoJZInBWKb9EgI4zLHpbQoeYcrsP+/X8/6ku5VSBkz7zHZeh1Ul8vwAKjYC5TbtM12fPMKlat
UOBMkl8axP7Ssgxx6IAAeY7uVL1h4jSbja9Sd6998Elj7YaOfTWSHl697BvbCBzGGzr4rLln2/sW
kkwg4Z5cK5btnqEohXMvHabrPwM+aBOf+RRj9mlgJ1izb8ZxAjMAMJDtnoPYpWPLr80GCDDa3ndw
VmDdBNCQFYiOx0YGgb/3T/L6ziyqpML4ZF0bx4U5ndcsMb/rJ6w/EGaOs9TzzrvgUrAQqlDJPOv7
QsATw7Zif9E4UnjS+R7YHvvIqx/gh8/fb27LUpf5Ys2vhaC+a6VJdxn1oWMgSNFBEGnrhmx5WY8/
HwK0c3g6kJ2I6gNPL87Y9WS2Io9wYbPTvlKBRRyTPRy9Pbj1K/MLITKdGhH8yrPsfqZR1jrazp4N
oorM8HEqgyravntSUoDvXuP+lvYWLx8zHCNcKy0BY5quoDTBzZcHPGZ7MK9I42xOK9Id/GG7TKwt
Qp+fGEw81/ef8KjE0WSYxBnpwtqRg3swL+xmfni6NzPxfx8Zasc3sucjDQSo+nHdmdHo7l0wLTjK
YNtY5J3u0LXoynNMSHMZhL3drANx1PkO1y4T8ij2PSWorDj2zkpMBBCWXnkiICdLkyMVRyV+XOTS
8rHlm7TZ//JNwiYu+FtYgGD7Y5lMbNPZizKUwJBckZur4e1n2J9EMSM116kT5YDcVaBSg36+ByQQ
aYTboUMpaKiT+ykl6qTqugDB+whudhTLrCURomwdICGPVzUP1OeIeKbURTn7hvXT71PzXMBGtA5e
jnd8haPVj3vfCOzS/xOeyM3CmkdqoXs+gSxR4QVbOQmuQsLw2QQ8OI8R5GaydoUJvnuKOiKdaBHn
7na6Le1jd9pdGOZHZaoATElUbMfCdEjd7LjaL8CE8+BSYZ2TLnpFFoHLj6S9HJKn7I97bn2doUoU
uH4Q3UWn4dO25Asza7+SuFIefBMwqiO0Sw/hFGZtY+OsJyV/rjiOSb2LXKmc7KRL6PebTEBiVnBy
sciU2HlndKN0CRHApiWuXtFaGAsiMiyie8R9Qxh7abuWmXuxWRCbPF3XT9XNgA2LcBvmyZKksUGO
AncgAeyWlrGhyq2osdIScRLp/8tH/+x5DBuoDUS1uF5zcLXl5iHWxVCM/cpAguUuLI9e84WNcIya
69n4UFCpGDi3gS+b4xAuGv1SNAjT4+rMkfUTWVQrZk30SXMWbvynfLUwdSs6dCcrpmqqT6cU0yrS
CGpIEHPXPRKhJ7t0hK8amE4Ol12TrNOkiCfychseRT9NEUmsOhtOIEWw+luFSDM1p4damaKJBMsQ
xEZlauRspDusliCK5vTDRr4mxR++oyPiPJBapIyuVT0y4srTsZfMUqYB3PICfQqSKr9ngJZNxVv1
C04UO0eYW1gJwHzmdFGcSCpyvvCU6yleWcal2tCeIauo8fi7AT+FakMR7Qv/UDhyEkYVoPXc6/M1
og1aUSg1hzuvnlrmUj64bze6d/WkBqJTzA8/s+bf5mWPl3iO8T8iAk7jaxX+4eh/Fxx7EbnGe6ZB
V9iXsm7mnncvrWh9wUz+TlLbSU/Ip4pgfU5OYT8+e48iLQCdXnz4GB6GO+YhcK7MWL549T4bQUBC
iBVHs+2zUVbyU4clf2YMRfrptMIG9J3x58jbKKrZP3ECztE0rZ2q2HA4YvIxIvP+DDo51YmkZE48
z1oZxdThMmpfnFnVZhRWmkEpDq6PGie2E/XzUJbq0btlnIaSe0nULkgow4SwmbRMixGwZi8zmE/o
gMTeASljOIrj3ZcWy/M7/7tjH2n89/v7SjeK8B6/traIyj8wBQaQbHuJqFeNAE/JqL1mj3QeXA+v
Uq2IfU1tn0j5+AtvLqUXyqXKqNHNWvf+1EtYCZeXdt5w0QaeW7V4UiE3RiMjnND/5r4JoazV8O7C
sqVWiy8EgfOPtAdVhma5cTskzhlXNSNeut1PFtO9mZsj+WX4YdtMpJmfGLlbkCMJcUBXOLdbb587
ynsKjzsAWfZZDo9K1/l3goR2rzqIg74jvthzY5cPDDCxpHc7Ewo4Um7FzZFv4NUOtxD0Zq0DwGGS
jsGonczH8gbjUyhpz1tfNa6WAE3pMSTJ1tpqAkGc0Hwnvw8JYKL7rhicHAcSrAys5c3UX+MMng/C
hO5V
`pragma protect end_protected
